package body Jtag2BSCANTbPkg is
  constant iSeq : TmsTdiArray := (
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"04000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"04000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffe2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffe3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000900", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"000000a9", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000040", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"ffa0a0a9", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000100", TDI => x"000000ff", nbits => 9),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000140", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"ffa0a0a9", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000100", TDI => x"000000ff", nbits => 9),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000240", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"ffa0a0a9", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000000", TDI => x"ffa0a0ff", nbits => 32),
( TMS => x"00000100", TDI => x"000000ff", nbits => 9),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000400", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"ffffffa9", nbits => 32),
( TMS => x"00000100", TDI => x"000000ff", nbits => 9),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000500", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"330000a9", nbits => 32),
( TMS => x"00000000", TDI => x"33000022", nbits => 32),
( TMS => x"00000000", TDI => x"33000022", nbits => 32),
( TMS => x"00000000", TDI => x"11001122", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"99889900", nbits => 32),
( TMS => x"00000000", TDI => x"88888888", nbits => 32),
( TMS => x"00000000", TDI => x"13021388", nbits => 32),
( TMS => x"00000000", TDI => x"99889902", nbits => 32),
( TMS => x"00000000", TDI => x"88888888", nbits => 32),
( TMS => x"00000000", TDI => x"13130288", nbits => 32),
( TMS => x"00000000", TDI => x"13130213", nbits => 32),
( TMS => x"00000000", TDI => x"13130213", nbits => 32),
( TMS => x"00000000", TDI => x"13130213", nbits => 32),
( TMS => x"00000000", TDI => x"bbbbaa13", nbits => 32),
( TMS => x"00000000", TDI => x"bbbbaabb", nbits => 32),
( TMS => x"00000000", TDI => x"bbbbbbbb", nbits => 32),
( TMS => x"00000000", TDI => x"bbbbbbbb", nbits => 32),
( TMS => x"00000000", TDI => x"000000bb", nbits => 32),
( TMS => x"00000000", TDI => x"00000080", nbits => 32),
( TMS => x"00000000", TDI => x"ffffff80", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"000002ff", nbits => 32),
( TMS => x"00000000", TDI => x"00000100", nbits => 32),
( TMS => x"00000000", TDI => x"ffffff00", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"000002ff", nbits => 32),
( TMS => x"00000000", TDI => x"00000100", nbits => 32),
( TMS => x"00000000", TDI => x"ffffff00", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"000000ff", nbits => 32),
( TMS => x"00000100", TDI => x"00000000", nbits => 9),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000800", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"000000a9", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000100", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00002000", TDI => x"00000000", nbits => 14),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"0000001f", TDI => x"00000000", nbits => 5 )
  );
  constant oSeq : TdoArray := (
( TDO => x"0000001f", nbits => 5),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"00000007", nbits => 3),
( TDO => x"0424a093", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00007fff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"08080fff", nbits => 32),
( TDO => x"81080738", nbits => 32),
( TDO => x"000000b0", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00007fff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"08080fff", nbits => 32),
( TDO => x"81080738", nbits => 32),
( TDO => x"000000b0", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"10080fff", nbits => 32),
( TDO => x"82080738", nbits => 32),
( TDO => x"ff805fb0", nbits => 32),
( TDO => x"21000001", nbits => 32),
( TDO => x"7fff8000", nbits => 32),
( TDO => x"801f8088", nbits => 32),
( TDO => x"001f8088", nbits => 32),
( TDO => x"f81f8089", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"10080fff", nbits => 32),
( TDO => x"82080738", nbits => 32),
( TDO => x"ff805fb0", nbits => 32),
( TDO => x"21000001", nbits => 32),
( TDO => x"7fff8000", nbits => 32),
( TDO => x"801f8088", nbits => 32),
( TDO => x"001f8088", nbits => 32),
( TDO => x"f81f8089", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"10080fff", nbits => 32),
( TDO => x"82080738", nbits => 32),
( TDO => x"ff805fb0", nbits => 32),
( TDO => x"21000001", nbits => 32),
( TDO => x"7fff8000", nbits => 32),
( TDO => x"801f8088", nbits => 32),
( TDO => x"001f8088", nbits => 32),
( TDO => x"f81f8089", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"000007ff", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00007fff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"08080fff", nbits => 32),
( TDO => x"81080738", nbits => 32),
( TDO => x"000000b0", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 32),
( TDO => x"00000000", nbits => 11),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000007ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00ffffff", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"000001ff", nbits => 9),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"000001ff", nbits => 9),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"000001ff", nbits => 9),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"000001ff", nbits => 9),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"ffffffff", nbits => 32),
( TDO => x"000001ff", nbits => 9),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"0001ffff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"00ffffff", nbits => 24),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"0000000f", nbits => 4),
( TDO => x"000003f1", nbits => 10),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"000187ff", nbits => 17),
( TDO => x"00000003", nbits => 2),
( TDO => x"00000007", nbits => 3),
( TDO => x"fff00fff", nbits => 32),
( TDO => x"000007ff", nbits => 32),
( TDO => x"00000800", nbits => 14),
( TDO => x"00000003", nbits => 2),
( TDO => x"0000001f", nbits => 5),
( TDO => x"00000001", nbits => 1),
( TDO => x"00000000", nbits => 5 )
  );
end package body Jtag2BSCANTbPkg;
