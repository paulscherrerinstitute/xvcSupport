package body Jtag2BSCANTbPkg is
  constant iSeq : TmsTdiArray := (
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"00000000", TDI => x"ffffffff", nbits => 32),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"04000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"00000000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"04000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffe2", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffc3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00800000", TDI => x"00000000", nbits => 24),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffff", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000003", TDI => x"00000000", nbits => 4),
( TMS => x"00000200", TDI => x"0000ffe3", nbits => 10),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00010000", TDI => x"0000f000", nbits => 17),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"00000001", TDI => x"00000000", nbits => 3),
( TMS => x"00000000", TDI => x"000000a9", nbits => 32),
( TMS => x"00000000", TDI => x"00000000", nbits => 32),
( TMS => x"00000400", TDI => x"00000000", nbits => 11),
( TMS => x"00000001", TDI => x"00000000", nbits => 2),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
( TMS => x"000000ff", TDI => x"00000000", nbits => 5),
( TMS => x"00000000", TDI => x"00000000", nbits => 1),
(TMS => x"0000001f", TDI => x"00000000", nbits => 5)
  );
end package body Jtag2BSCANTbPkg;
